module Forward_ALU_Mux
(
  input [31:0] reg_ex_in,
  input [31:0] reg_wb_in,
  input [31:0] reg_mem_in,
  input [1:0] forward_control_in,
  output reg [31:0] reg_out
);
	always @(*) begin
		case (forward_control_in)
        2'b01 : reg_out <= reg_wb_in;
        2'b10 : reg_out <= reg_mem_in;
        default : reg_out <= reg_ex_in;
      endcase
	end
endmodule